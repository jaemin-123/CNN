`timescale 1ns / 1ps

module requantizer #(
    parameter IN_W = 24,
    parameter OUT_W = 8,
    parameter MULTIPLIER = 350896, // ���� �� ���� (Top���� ��������� �����ϰ�)
    parameter SHIFT = 16
)(
    input  wire clk, rst_n, valid_in,
    input  wire signed [IN_W-1:0] data_in,
    
    output reg  valid_out,
    output reg  signed [OUT_W-1:0] data_out
);

    // ============================================================
    // [Stage 1] �Է� �������� (Routing Delay ����)
    // ============================================================
    reg signed [IN_W-1:0] r_data_in;
    reg r_valid_in;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            r_data_in  <= 0;
            r_valid_in <= 0;
        end else begin
            r_data_in  <= data_in;
            r_valid_in <= valid_in;
        end
    end

    // ============================================================
    // [Stage 2] ���� �������� (Logic Delay�� �ٽ� - DSP ��� ���)
    // ============================================================
    reg signed [63:0] r_mult_res; // ���� ����� �˳��ϰ� 64��Ʈ
    reg r_valid_mult;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            r_mult_res   <= 0;
            r_valid_mult <= 0;
        end else begin
            if (r_valid_in) begin
                // ���⼭ ������ �����̰� �߻��ϴ� ������ �����ϰ� ����
                r_mult_res   <= r_data_in * $signed(MULTIPLIER);
                r_valid_mult <= 1;
            end else begin
                r_mult_res   <= 0;
                r_valid_mult <= 0;
            end
        end
    end

    // ============================================================
    // [Combinational Logic] �ݿø� & ����Ʈ & Ŭ���� (��길 ��)
    // ============================================================
    wire signed [63:0] rounded;
    wire signed [63:0] shifted;
    reg  signed [OUT_W-1:0] clamped_val; // ���� ���� �� (���� �������� �ƴ�)

    // 1. �ݿø� (����ڴ� ���� �ڵ� ����)
    generate
        if (SHIFT > 0) begin : GEN_ROUND
            assign rounded = r_mult_res + (1 << (SHIFT - 1));
        end else begin : GEN_NO_ROUND
            assign rounded = r_mult_res;
        end
    endgenerate

    // 2. ����Ʈ
    assign shifted = rounded >>> SHIFT;

    // 3. Ŭ���� (Saturate) - ���� ȸ�η� ����
    always @(*) begin
        if (shifted > 127)      
            clamped_val = 8'sd127;
        else if (shifted < -128) 
            clamped_val = -8'sd128;
        else                     
            clamped_val = shifted[OUT_W-1:0];
    end

    // ============================================================
    // [Stage 3] ��� �������� (���� ��� ��������)
    // ============================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            data_out  <= 0;
            valid_out <= 0;
        end else begin
            // ���� Ŭ���� ���� �������Ϳ� ��Ƽ� ��� (Ÿ�̹� Ȯ��)
            if (r_valid_mult) begin
                data_out  <= clamped_val;
                valid_out <= 1;
            end else begin
                data_out  <= 0;
                valid_out <= 0;
            end
        end
    end

endmodule