`timescale 1ns / 1ps

module cnn_multichannel_top #(
    parameter DATA_W = 8,
    parameter ACC_W  = 24,
    parameter IMG_W  = 28
)(
    input  wire clk, rst_n, valid_in,
    input  wire [DATA_W-1:0] data_in,
    
    output wire fc_done,
    output wire [3:0] final_digit
    
    // (������)
//    output wire signed [DATA_W-1:0] l2_ch0_out, l2_ch1_out, l2_ch2_out,
//    output wire l2_valid_out
);

    // ====================================================================
    // Bias (No-Bias Model)
    // ====================================================================
    wire signed [23:0] l1_bias [0:2];
    assign l1_bias[0] = 0; assign l1_bias[1] = 0; assign l1_bias[2] = 0;

    wire signed [23:0] l2_bias [0:2];
    assign l2_bias[0] = 0; assign l2_bias[1] = 0; assign l2_bias[2] = 0;
    
    // ====================================================================
    // �� [����] ���� ROM ���� (�ܺ� �Է� ��� ���)
    // ====================================================================
//    reg  [9:0] rom_addr;
//    wire signed [7:0] rom_data;
    
//    // �̹��� ROM �ν��Ͻ�
//    single_image_rom u_test_rom (
//        .clk(clk),
//        .addr(rom_addr),
//        .data_out(rom_data)
//    );

//    reg signed [DATA_W-1:0] internal_data;
//    reg internal_valid;
    
//    // �����͸� �о�ͼ� CNN���� �־��ִ� ������ ���� �ӽ�
//    reg [1:0] state;
    
//    always @(posedge clk or negedge rst_n) begin
//        if (!rst_n) begin
//            rom_addr <= 0;
//            state <= 0;
//            internal_valid <= 0;
//            internal_data <= 0;
//        end else begin
//            case(state)
//                0: begin // ��� ����
//                    internal_valid <= 0;
//                    rom_addr <= 0;
//                    if (valid_in) state <= 1; // ��ư ������ ����
//                end
                
//                1: begin // �б� ����
//                    internal_data <= rom_data; // ROM ������ -> CNN �Է�
//                    internal_valid <= 1;       // Valid ��ȣ ON
                    
//                    if (rom_addr < 783) begin
//                        rom_addr <= rom_addr + 1;
//                    end else begin
//                        state <= 0; // 784�� �� �־����� ��
//                    end
//                end
//            endcase
//        end
//    end
    
    // ====================================================================
    // 0. Pre-processing Unit (��ó�� ��� �߰�)
    // ====================================================================
    wire pre_valid;
    wire signed [DATA_W-1:0] pre_data;
    
    preprocessing_unit u_pre (
        .clk(clk),
        .rst_n(rst_n),
        .valid_in(valid_in),
        .raw_data_in(data_in),
        .valid_out(pre_valid),
        .data_out(pre_data)
    );

    // ====================================================================
    // ���� ���� ���� (�Է��� pre_valid, pre_data�� ����)
    // ====================================================================
    
    // Input Buffer
    reg signed [DATA_W-1:0] internal_data;
    reg internal_valid;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            internal_valid <= 0;
            internal_data  <= 0;
        end else begin
            // �� ������: �ܺ� �Է� ��� ��ó�� ��� ����� ����
            internal_valid <= pre_valid;
            internal_data  <= pre_data; 
        end
    end
    
    // Weight ROM
    wire [DATA_W*75-1:0]  l1_w_flat;
    wire [DATA_W*225-1:0] l2_w_flat;
    wire [DATA_W*480-1:0] fc_w_flat; 
    
    weight_rom #(.DATA_W(DATA_W)) w_rom (
        .l1_weights_flat(l1_w_flat),
        .l2_weights_flat(l2_w_flat),
        .fc_weights_flat(fc_w_flat)
    );

    // Layer 1
    wire [DATA_W*25-1:0] l1_win_flat;
    wire l1_win_valid;
    
    line_buffer_wrapper_5x5 #(.W(IMG_W), .D(DATA_W)) lb_l1 (
        .clk(clk), .rst_n(rst_n), 
        .d_in(internal_data), .v_in(internal_valid),  
        .win_flat_vec(l1_win_flat), .v_out(l1_win_valid)
    );

    wire signed [DATA_W-1:0] l1_pool_out[0:2];
    wire l1_pool_valid[0:2];

    genvar i;
    generate
        for (i=0; i<3; i=i+1) begin : GEN_L1
            wire signed [ACC_W-1:0] conv_y;
            wire conv_valid;
            
            wire signed [DATA_W-1:0] w[0:24];
            wire signed [DATA_W-1:0] k[0:24];
            genvar j;
            for(j=0; j<25; j=j+1) begin : ASSIGN_L1
                assign w[j] = l1_win_flat[(25-j)*DATA_W-1 -: DATA_W];
                assign k[j] = l1_w_flat[ (75 - i*25 - j)*DATA_W - 1 -: DATA_W ];
            end
            
            conv5x5_single_filter #(.DATA_BITS(DATA_W), .SUM_BITS(ACC_W)) conv_inst (
                .clk(clk), .rst_n(rst_n), .valid_in(l1_win_valid),
                .p00(w[0]), .p01(w[1]), .p02(w[2]), .p03(w[3]), .p04(w[4]),
                .p10(w[5]), .p11(w[6]), .p12(w[7]), .p13(w[8]), .p14(w[9]),
                .p20(w[10]),.p21(w[11]),.p22(w[12]),.p23(w[13]),.p24(w[14]),
                .p30(w[15]),.p31(w[16]),.p32(w[17]),.p33(w[18]),.p34(w[19]),
                .p40(w[20]),.p41(w[21]),.p42(w[22]),.p43(w[23]),.p44(w[24]),
                .k00(k[0]), .k01(k[1]), .k02(k[2]), .k03(k[3]), .k04(k[4]),
                .k10(k[5]), .k11(k[6]), .k12(k[7]), .k13(k[8]), .k14(k[9]),
                .k20(k[10]),.k21(k[11]),.k22(k[12]),.k23(k[13]),.k24(k[14]),
                .k30(k[15]),.k31(k[16]),.k32(k[17]),.k33(k[18]),.k34(k[19]),
                .k40(k[20]),.k41(k[21]),.k42(k[22]),.k43(k[23]),.k44(k[24]),
                .bias(l1_bias[i]),
                .valid_out(conv_valid), .y(conv_y)
            );

            wire rq_valid_out;
            wire signed [DATA_W-1:0] rq_y;
            requantizer #(.IN_W(ACC_W), .OUT_W(DATA_W), .MULTIPLIER(59), .SHIFT(16)) rq (
                .clk(clk), .rst_n(rst_n), 
                .valid_in(conv_valid), .data_in(conv_y), 
                .valid_out(rq_valid_out), .data_out(rq_y)
            );

            wire signed [DATA_W-1:0] relu_y;
            wire relu_valid;
            relu #(.DATA_W(DATA_W)) relu_block (
                .clk(clk), .rst_n(rst_n), 
                .valid_in(rq_valid_out), .in(rq_y),
                .valid_out(relu_valid), .out(relu_y)
            );

            wire signed [DATA_W-1:0] mp_p00, mp_p01, mp_p10, mp_p11;
            wire mp_valid_in;
            line_buffer_2x2 #(.DATA_BITS(DATA_W), .DATA_W(24)) lb2 (
                .clk(clk), .rst_n(rst_n), .data_in(relu_y), .valid_in(relu_valid),
                .p00(mp_p00), .p01(mp_p01), .p10(mp_p10), .p11(mp_p11), .window_valid(mp_valid_in)
            );
            maxpool2x2_core #(.DATA_W(DATA_W)) mp (
                .clk(clk), .rst_n(rst_n), .valid_in(mp_valid_in),
                .p00(mp_p00), .p01(mp_p01), .p10(mp_p10), .p11(mp_p11),
                .valid_out(l1_pool_valid[i]), .y(l1_pool_out[i])
            );
        end
    endgenerate

    // Layer 2
    wire [DATA_W*25-1:0] l2_win_flat_ch0, l2_win_flat_ch1, l2_win_flat_ch2;
    wire l2_v0, l2_v1, l2_v2;
    wire l2_common_valid = l2_v0 & l2_v1 & l2_v2;

    line_buffer_wrapper_5x5 #(.W(12), .D(DATA_W)) lb_l2_c0 (
        .clk(clk), .rst_n(rst_n), .d_in(l1_pool_out[0]), .v_in(l1_pool_valid[0]), 
        .win_flat_vec(l2_win_flat_ch0), .v_out(l2_v0)
    );
    line_buffer_wrapper_5x5 #(.W(12), .D(DATA_W)) lb_l2_c1 (
        .clk(clk), .rst_n(rst_n), .d_in(l1_pool_out[1]), .v_in(l1_pool_valid[1]), 
        .win_flat_vec(l2_win_flat_ch1), .v_out(l2_v1)
    );
    line_buffer_wrapper_5x5 #(.W(12), .D(DATA_W)) lb_l2_c2 (
        .clk(clk), .rst_n(rst_n), .d_in(l1_pool_out[2]), .v_in(l1_pool_valid[2]), 
        .win_flat_vec(l2_win_flat_ch2), .v_out(l2_v2)
    );

    wire signed [DATA_W-1:0] l2_res[0:2];
    wire l2_res_valid[0:2];
    
    // =========================================================
    // [DEBUG] Layer 2 Input Window Monitor (Ch0�� Ȯ��)
    // =========================================================
    // Layer 2�� ù ��° ������ ����� ��, 5x5 ������ ���� ���ϴ�.
    
//    always @(posedge clk) begin
//        // l2_common_valid�� 1�� �Ǵ� ������ ���� �������Դϴ�.
//        if (l2_common_valid) begin
//            // �ʹ� ���� ������ ���� ����ϱ� ó�� 3���� ����ϴ�.
//            if ($time < 50000) begin // ������ �ð� ����
//                 $display("\n[Verilog L2 Input Window Ch0]");
//                 // 5x5 ������� l2_win_flat_ch0�� ��źȭ�Ǿ� �ֽ��ϴ�.
//                 // ���� �ֱ� ��(Row4, Col4)���� �������� ������� �� ������ Ȯ�� �ʿ�
//                 // ���⼭�� 5x5 �� ���� �߽ɰ�(Center)�̳� ù ��° ���� ���ô�.
                 
//                 // l2_win_flat_ch0 ����: [p00, p01... p44] �������� Ȯ��
//                 // ���� Line Buffer Wrapper���� ����� �� Flatten �մϴ�.
                 
//                 $display("Window Flat: %h", l2_win_flat_ch0);
//            end
//        end
//    end

    generate
        for (i=0; i<3; i=i+1) begin : GEN_L2
            wire signed [ACC_W-1:0] sum_y;
            wire sum_valid;
            
            wire [DATA_W*75-1:0] current_ch_weights;
            assign current_ch_weights = l2_w_flat[ (225 - i*75)*DATA_W - 1 -: DATA_W*75 ];
//            assign current_ch_weights = l2_w_flat[ (i*75)*DATA_W +: DATA_W*75 ];
            
            conv_3ch_sum_PE #(.DATA_W(DATA_W), .ACC_W(ACC_W)) pe_inst (
                .clk(clk), .rst_n(rst_n), .valid_in(l2_common_valid),
                .ch0_flat(l2_win_flat_ch0),
                .ch1_flat(l2_win_flat_ch1),
                .ch2_flat(l2_win_flat_ch2),
                .weights_flat(current_ch_weights),
                .sum_out(sum_y), .valid_out(sum_valid)
            );
            // �ڡڡ� [DEBUG] ���Ⱑ �ٽ��Դϴ�! �ڡڡ�
            // i==0 (ù��° ��� ä��)�� ����� ���ϴ�.
//            always @(posedge clk) begin
//                if (i == 0 && sum_valid) begin
//                    // �ʹ� ���� ������ ���� ����ϱ� �ʹ� 10����
//                    if ($time < 500000) 
//                        $display("[Verilog L2 Raw] Val: %d", $signed(sum_y));
//                end
//            end
            
            wire signed [ACC_W-1:0] sum_y_biased;
            assign sum_y_biased = sum_y + l2_bias[i];

            wire rq_valid_l2;
            wire signed [DATA_W-1:0] rq_y;
            
            requantizer #(.IN_W(ACC_W), .OUT_W(DATA_W), .MULTIPLIER(97), .SHIFT(16)) rq_l2 (
                .clk(clk), .rst_n(rst_n), 
                .valid_in(sum_valid), .data_in(sum_y_biased),
                .valid_out(rq_valid_l2), .data_out(rq_y)
            );
            
//            always @(posedge clk) begin
//                // rq_valid_l2�� �� ������ ��� ä�ο��� ���� ���� �������� Ȯ��
//                if (rq_valid_l2) begin
//                    $display("[Verilog L2 Check] Ch %0d | Val: %d", i, $signed(rq_y));
//                end
//            end
            
            // �ڡڡ� [DEBUG] Requantizer ��� Ȯ�� (������) �ڡڡ�
//            always @(posedge clk) begin
//                if (i == 0 && rq_valid_l2) begin
//                    // ������ 64�� ������ Ȯ��
//                    if ($time < 500000) 
//                        $display("[Verilog L2 Requant] Val: %d", $signed(rq_y));
//                end
//            end

            wire signed [DATA_W-1:0] relu_y;
            wire relu_valid;
            relu #(.DATA_W(DATA_W)) relu_block_l2 (
                .clk(clk), .rst_n(rst_n), 
                .valid_in(rq_valid_l2), .in(rq_y),
                .valid_out(relu_valid), .out(relu_y)
            );
            
            // �ڡڡ� [DEBUG] ReLU ��� Ȯ�� (Ch0��) �ڡڡ�
//            always @(posedge clk) begin
//                if (i == 0 && relu_valid) begin
//                    if ($time < 500000) 
//                        $display("[Verilog L2 ReLU] Val: %d", $signed(relu_y));
//                end
//            end

            wire signed [DATA_W-1:0] mp_p00, mp_p01, mp_p10, mp_p11;
            wire mp_v;
            line_buffer_2x2 #(.DATA_BITS(DATA_W), .DATA_W(8)) lb2_l2 (
                .clk(clk), .rst_n(rst_n), .data_in(relu_y), .valid_in(relu_valid),
                .p00(mp_p00), .p01(mp_p01), .p10(mp_p10), .p11(mp_p11), .window_valid(mp_v)
            );
            maxpool2x2_core #(.DATA_W(DATA_W)) mp_l2 (
                .clk(clk), .rst_n(rst_n), .valid_in(mp_v),
                .p00(mp_p00), .p01(mp_p01), .p10(mp_p10), .p11(mp_p11),
                .valid_out(l2_res_valid[i]), .y(l2_res[i])
            );
//            always @(posedge clk) begin
//                if (i == 0) begin
//                    if (sum_valid)    $display("[L2_DEBUG] RAW_SUM: %d", $signed(sum_y));
//                    if (rq_valid_l2)  $display("[L2_DEBUG] REQUANT: %d", $signed(rq_y));
//                    if (relu_valid)   $display("[L2_DEBUG] RELU   : %d", $signed(relu_y));
//                    if (l2_res_valid[0]) $display("[L2_DEBUG] MAXPOOL: %d <--- FC �Ա�", $signed(l2_res[0]));
//                end
//            end
        end
    endgenerate
    
    // ====================================================================
    // FC Layer (Final)
    // ====================================================================
    wire signed [DATA_W-1:0] fc_raw_data;
    wire fc_raw_valid;
    
    // ====================================================================
    // �� [DEBUG] P2S �Է� 3ä�� ���� ���� ��
    // ====================================================================
    
//    always @(posedge clk) begin
//        // 3�� �� �ϳ��� ��ȿ�ϸ� ���ϴ�.
//        if (l2_res_valid[0] || l2_res_valid[1] || l2_res_valid[2]) begin
//             $display("[P2S INPUT Check] Ch0: %d | Ch1: %d | Ch2: %d", 
//                      $signed(l2_res[0]), $signed(l2_res[1]), $signed(l2_res[2]));
//        end
//    end
    
    // 1. Parallel to Serial (�ܼ� ����)
    parallel_to_serial #(.DATA_W(DATA_W)) u_serializer (
        .clk(clk), .rst_n(rst_n),
        .din_0(l2_res[0]), .vin_0(l2_res_valid[0]),
        .din_1(l2_res[1]), .vin_1(l2_res_valid[1]),
        .din_2(l2_res[2]), .vin_2(l2_res_valid[2]),
        .dout(fc_raw_data), .vout(fc_raw_valid)
    );
    
    // �ڡڡ� [DEBUG] MaxPool ��� (P2S �Է�) Ȯ�� �ڡڡ�
    // 58(����)���� 85(������)���� Ȯ���ϴ� ������ �ڵ�
//    always @(posedge clk) begin
//        // l2_res_valid[0]�� MaxPool�� ��ȿ�� �����͸� ���� �� 1�� �˴ϴ�.
//        if (l2_res_valid[0]) begin
//             $display("[Verilog MaxPool Out] Ch0 Val: %d", $signed(l2_res[0]));
//        end
//    end

    // �ڡڡ� [FINAL CHECK] FC �Է� ������ ���� �ڡڡ�
    // P2S�� ����ؼ� FC�� ���� ���� ������
//    reg [31:0] check_cnt;
//    always @(posedge clk or negedge rst_n) begin
//        if(!rst_n) check_cnt <= 0;
//        else if(fc_raw_valid) begin
//            $display("[Verilog FC Input] Index %0d: %d", check_cnt, $signed(fc_raw_data));
//            check_cnt <= check_cnt + 1;
//        end
//    end

    // �ڡڡ� [�ٽ�] 48�� ī���� & ����Ʈ (Safety Gate) �ڡڡ�
    // ������ �����Ͱ� ������ ���� ���� ���� 0~47�������� ���� �����ݴϴ�.
    
    reg [5:0] fc_input_cnt;
//    reg fc_gated_valid;
//    reg signed [DATA_W-1:0] fc_gated_data; // �� ������ ����ȭ�� �������� �߰�
    
    wire fc_gated_valid;
    wire signed [DATA_W-1:0] fc_gated_data; // �� ������ ����ȭ�� �������� �߰�

//    always @(posedge clk or negedge rst_n) begin
//        if (!rst_n) begin
//            fc_input_cnt <= 0;
//            fc_gated_valid <= 0;
//            fc_gated_data <= 0; // ���� �߰�
//        end else begin
//            if (fc_raw_valid && fc_input_cnt < 48) begin
//                fc_gated_valid <= 1;
//                fc_gated_data  <= fc_raw_data; // �� �����͵� ���⼭ ĸó (1Ŭ�� ������)
//                fc_input_cnt   <= fc_input_cnt + 1;
//            end else begin
//                fc_gated_valid <= 0;
//                fc_gated_data  <= 0; // (���û���) �����ϰ� 0 ó��
//            end
//        end
//    end
    assign fc_gated_valid = fc_raw_valid; 
    assign fc_gated_data  = fc_raw_data;

    // 2. FC Layer ���� ����
    fc_layer #(.DATA_W(DATA_W), .MULTIPLIER(346)) fc_inst (
        .clk(clk),
        .rst_n(rst_n),
        .valid_in(fc_gated_valid), 
        .data_in(fc_gated_data),     // �� fc_raw_data ��� fc_gated_data ����
        .weights_flat(fc_w_flat), 
        .valid_out(fc_done),
        .predicted_class(final_digit)
    );
    
    // ====================================================================
    // �� [DEBUG] ���̽� �񱳿� ������ ���� (�ڵ� ī���� �߰�)
    // ====================================================================
//    integer f;
//    integer dbg_img_cnt; // ���ο��� �̹��� ������ ���� ���� ����

//    initial begin
//        f = $fopen("verilog_fc_input_dump.txt", "w");
//        dbg_img_cnt = 0;
//    end

//    always @(posedge clk) begin
//        // fc_gated_valid�� 1�� �� (FC�� �����Ͱ� ���� ����)
//        if (fc_gated_valid) begin
//            // ���Ͽ� ���: �̹�����ȣ, �ε���(0~47), ��
//            // �� �߿�: fc_raw_data�� �ƴ϶� Ÿ�̹� ���� 'fc_gated_data'�� ���� �մϴ�.
//            $fwrite(f, "Img_%0d, Idx_%0d, Val_%d\n", dbg_img_cnt, fc_input_cnt, $signed(fc_gated_data));

//            // ���� ������ 47�� �ε������ٸ�, �̹��� ī��Ʈ ����
//            if (fc_input_cnt == 47) begin
//                dbg_img_cnt = dbg_img_cnt + 1;
//                $fwrite(f, "--------------------------------\n"); // ���м�
//            end
//        end
//    end

endmodule