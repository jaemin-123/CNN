`timescale 1ns / 1ps

module single_image_rom (
    input wire clk,
    input wire [9:0] addr,  // 0~783 (784�� �ȼ�)
    output reg signed [7:0] data_out
);
    // 1�� �̹��� (784����Ʈ) ���� ����
    reg [7:0] memory [0:783];

    initial begin
        // �� �߿�: ���� ��� hex ���� �� �ϳ��� �����ؼ� "image_1.hex"�� ���弼��
        // Ȥ�� ���� hex ������ �״�� ����, ó�� 784�ٸ� �����ϴ�.
        $readmemh("D:/01_work_verilog/01_CNN/images_100.hex", memory);
    end

    always @(posedge clk) begin
        data_out <= memory[addr];
    end
endmodule