`timescale 1ns / 1ps

module weight_rom #(
    parameter DATA_W = 8
)(
    output wire [DATA_W*75-1:0] l1_weights_flat,
    output wire [DATA_W*225-1:0] l2_weights_flat
);

    reg [DATA_W*75-1:0]  l1_storage;
    reg [DATA_W*225-1:0] l2_storage;

    assign l1_weights_flat = l1_storage;
    assign l2_weights_flat = l2_storage;

    initial begin
        // =================================================================
        // [1] Layer 1 Weights (�� 75��) - C ���� �� ����
        // =================================================================
        l1_storage = {
            // Filter 0 (Index 0~24)
             8'sd7,  8'sd76,  8'sd93,  8'sd63,  8'sd18, 
            -8'sd23, 8'sd109, 8'sd40,  8'sd100, -8'sd37, 
             8'sd74, 8'sd49,  8'sd108, 8'sd55,  8'sd70, 
             8'sd73, 8'sd127, 8'sd74,  8'sd47,  8'sd28, 
             8'sd113,8'sd120, 8'sd44,  8'sd15, -8'sd10,

            // Filter 1 (Index 25~49)
            -8'sd68, -8'sd32,  8'sd44,  8'sd127, 8'sd86, 
            -8'sd10, -8'sd32,  8'sd14,  8'sd47,  8'sd107, 
            -8'sd101,-8'sd46, -8'sd27, -8'sd5,   8'sd66, 
            -8'sd89, -8'sd117,-8'sd39,  8'sd15,  8'sd50, 
            -8'sd31, -8'sd40, -8'sd90, -8'sd50,  8'sd19,

            // Filter 2 (Index 50~74)
             8'sd105, 8'sd127, 8'sd78,  8'sd30, -8'sd39, 
             8'sd21,  8'sd59,  8'sd116, 8'sd102,-8'sd24, 
            -8'sd18,  8'sd20,  8'sd32,  8'sd76,  8'sd11, 
            -8'sd99, -8'sd73, -8'sd40,  8'sd34,  8'sd63, 
            -8'sd65, -8'sd53, -8'sd44, -8'sd19,  8'sd80
        };

        // =================================================================
        // [2] Layer 2 Weights (�� 225��) - C ���� �� ����
        // =================================================================
        l2_storage = {
            // -----------------------------------------------------------
            // Output Channel 0 (�� 75��)
            // -----------------------------------------------------------
             8'sd1,  -8'sd16,  8'sd3,  -8'sd15, -8'sd33, 
             8'sd4,  -8'sd25, -8'sd23, -8'sd41, -8'sd62, 
            -8'sd14,  8'sd5,  -8'sd3,   8'sd21, -8'sd30, 
            -8'sd48, -8'sd28,  8'sd5,   8'sd21,  8'sd12, 
             8'sd27,  8'sd19,  8'sd9,   8'sd2,  -8'sd8, 
            -8'sd14, -8'sd23, -8'sd78, -8'sd87, -8'sd38, 
            -8'sd19, -8'sd43, -8'sd36, -8'sd1,   8'sd51, 
            -8'sd13,  8'sd5,   8'sd38,  8'sd59, -8'sd63, 
             8'sd27,  8'sd48,  8'sd29,  8'sd54,  8'sd0, 
             8'sd3,  -8'sd17, -8'sd6,  -8'sd19,  8'sd14, 
             8'sd28, -8'sd17, -8'sd8,   8'sd15,  8'sd55, 
             8'sd33,  8'sd31,  8'sd39,  8'sd89,  8'sd75, 
            -8'sd2,   8'sd56,  8'sd65,  8'sd127, 8'sd70, 
             8'sd13,  8'sd87,  8'sd97,  8'sd62,  8'sd39, 
             8'sd28,  8'sd20,  8'sd38,  8'sd16,  8'sd25,

            // -----------------------------------------------------------
            // Output Channel 1 (�� 75��)
            // -----------------------------------------------------------
            -8'sd43,  8'sd38,  8'sd37,  8'sd38,  8'sd43, 
             8'sd47,  8'sd17,  8'sd41,  8'sd18,  8'sd39, 
             8'sd10,  8'sd14,  8'sd3,  -8'sd43, -8'sd56, 
             8'sd5,  -8'sd14, -8'sd27, -8'sd31, -8'sd37, 
            -8'sd50, -8'sd22, -8'sd31,  8'sd2,  -8'sd3, 
             8'sd17,  8'sd14,  8'sd11, -8'sd57, -8'sd127,
             8'sd28,  8'sd37,  8'sd33,  8'sd74,  8'sd104,
             8'sd14,  8'sd41,  8'sd54,  8'sd26,  8'sd17, 
             8'sd37,  8'sd19,  8'sd13, -8'sd56, -8'sd78, 
             8'sd8,   8'sd14,  8'sd15, -8'sd22, -8'sd42, 
            -8'sd29, -8'sd26, -8'sd26, -8'sd49, -8'sd54, 
             8'sd31,  8'sd9,  -8'sd2,  -8'sd7,   8'sd42, 
             8'sd15,  8'sd19,  8'sd1,   8'sd28,  8'sd23, 
             8'sd60,  8'sd16, -8'sd31, -8'sd5,  -8'sd9, 
            -8'sd26, -8'sd8,  -8'sd44, -8'sd12, -8'sd7,

            // -----------------------------------------------------------
            // Output Channel 2 (�� 75��)
            // -----------------------------------------------------------
             8'sd10,  8'sd106, 8'sd127, 8'sd46,  8'sd8, 
             8'sd92,  8'sd101,-8'sd13, -8'sd40, -8'sd9, 
             8'sd15,  8'sd2,  -8'sd64, -8'sd38, -8'sd4, 
             8'sd34,  8'sd14, -8'sd9,  -8'sd5,  -8'sd25, 
             8'sd41,  8'sd54,  8'sd40,  8'sd16, -8'sd59, 
             8'sd40, -8'sd16, -8'sd61, -8'sd96, -8'sd48, 
             8'sd49, -8'sd60, -8'sd82, -8'sd12,  8'sd44, 
             8'sd72, -8'sd71,  8'sd11,  8'sd79,  8'sd48, 
             8'sd40,  8'sd110,-8'sd5,   8'sd89,  8'sd47, 
             8'sd61,  8'sd62,  8'sd15, -8'sd3,   8'sd20, 
            -8'sd52, -8'sd104,-8'sd32,  8'sd28,  8'sd28, 
            -8'sd48, -8'sd118, 8'sd10, -8'sd22, -8'sd34, 
            -8'sd38, -8'sd86, -8'sd85, -8'sd34, -8'sd6, 
            -8'sd11, -8'sd10, -8'sd22, -8'sd73,  8'sd21, 
             8'sd27, -8'sd3,   8'sd10, -8'sd37, -8'sd38
        };
    end
endmodule