//`timescale 1ns / 1ps

//module tb_cnn_1000;

//    // ==========================================
//    // Parameters
//    // ==========================================
//    parameter DATA_W = 8;
//    parameter IMG_W  = 28;
//    parameter CLK_PERIOD = 8;
    
//    // �� ������: 1000�� �׽�Ʈ
//    parameter NUM_TEST = 1000; 

//    reg clk, rst_n, valid_in;
//    reg signed [DATA_W-1:0] data_in;
//    wire fc_done;
//    wire [3:0] final_digit;

//    // DUT ����
//    cnn_multichannel_top #(.DATA_W(DATA_W), .IMG_W(IMG_W)) dut (
//        .clk(clk), .rst_n(rst_n), .valid_in(valid_in), .data_in(data_in),
//        .fc_done(fc_done), .final_digit(final_digit)
//    );

//    // �� ������: �޸� ũ�� ���� (784 * 1000)
//    reg [DATA_W-1:0] all_images [0 : 784*1000 - 1];
//    reg [7:0]        all_labels [0 : 999];

//    // Clock Generation
//    initial clk = 0;
//    always #(CLK_PERIOD/2) clk = ~clk;

//    integer img_idx, px_idx;
//    integer correct_cnt;
//    integer base_addr;
//    reg [3:0] correct_label;

//    initial begin
//        // �� ���ϸ� Ȯ�� (��δ� �ùķ��̼� ȯ�濡 �����ּ���)
//        $readmemh("raw_images_1000.hex", all_images);
//        $readmemh("labels_1000.hex", all_labels);
        
//        // �ʱ�ȭ
//        rst_n = 0; valid_in = 0; data_in = 0;
//        correct_cnt = 0;

//        #100; rst_n = 1; #20;

//        $display("\n========================================");
//        $display(" Start Testing %0d Images...", NUM_TEST);
//        $display("========================================\n");

//        for (img_idx = 0; img_idx < NUM_TEST; img_idx = img_idx + 1) begin
            
//            // �̹��� �ٲ� ������ ���� (�����ϰ�)
//            rst_n = 0; #20; rst_n = 1; #20;

//            correct_label = all_labels[img_idx][3:0];
//            base_addr = img_idx * 784;

//            // �ȼ� ����
//            for (px_idx = 0; px_idx < 784; px_idx = px_idx + 1) begin
//                @(negedge clk);
//                valid_in = 1;
//                data_in = all_images[base_addr + px_idx];
//            end

//            @(negedge clk);
//            valid_in = 0;
//            data_in = 0;

//            // ��� ���
//            wait(fc_done);
//            @(posedge clk);

//            // ä��
//            if (final_digit == correct_label) begin
//                correct_cnt = correct_cnt + 1;
//            end else begin
//                // Ʋ�� ��� ���
//                $display("Img %0d: FAIL (Pred: %d, True: %d)", img_idx, final_digit, correct_label);
//            end
            
//            // ���� ��Ȳ ��� (100������)
//            if ((img_idx + 1) % 100 == 0) begin
//                $display("Process: %0d / %0d done... (Current Acc: %0d %%)", 
//                         img_idx + 1, NUM_TEST, correct_cnt * 100 / (img_idx + 1));
//            end

//            #200; // ���� �̹��� �� ������
//        end

//        $display("\n========================================");
//        $display(" Test Finished!");
//        $display(" Total Images: %0d", NUM_TEST);
//        $display(" Correct:      %0d", correct_cnt);
//        // �Ҽ��� ����� �� �Ǵ� ���������� �뷫 ���
//        $display(" Accuracy:      %0d.%0d %%", (correct_cnt * 100 / NUM_TEST), (correct_cnt * 1000 / NUM_TEST) % 10);
//        $display("========================================");
        
//        $finish;
//    end

//endmodule

`timescale 1ns / 1ps

module tb_cnn_10000; // ��� �̸��� 10000���� �����ϸ� ������ �����ϴ�

    // ==========================================
    // Parameters
    // ==========================================
    parameter DATA_W = 8;
    parameter IMG_W  = 28;
    parameter CLK_PERIOD = 8;
    
    // �� 10,000�� �׽�Ʈ ����
    parameter NUM_TEST = 10000; 

    reg clk, rst_n, valid_in;
    reg signed [DATA_W-1:0] data_in;
    wire fc_done;
    wire [3:0] final_digit;

    // DUT ����
    cnn_multichannel_top #(.DATA_W(DATA_W), .IMG_W(IMG_W)) dut (
        .clk(clk), .rst_n(rst_n), .valid_in(valid_in), .data_in(data_in),
        .fc_done(fc_done), .final_digit(final_digit)
    );

    // ==========================================
    // �� [�߿�] �޸� ũ�� ���� (10,000�� �з� Ȯ��)
    // ==========================================
    // 784�ȼ� * 10,000�� = 7,840,000�� �ּ� �ʿ�
    reg [DATA_W-1:0] all_images [0 : 784*10000 - 1]; 
    
    // ���� �� 10,000��
    reg [7:0]        all_labels [0 : 9999];

    // Clock Generation
    initial clk = 0;
    always #(CLK_PERIOD/2) clk = ~clk;

    integer img_idx, px_idx;
    integer correct_cnt;
    integer base_addr;
    reg [3:0] correct_label;

    initial begin
        // ���� �ε� (���ε����ֽ� ���ϸ�� ��ġ)
        $display("Loading Hex Files...");
        $readmemh("raw_images_10000.hex", all_images);
        $readmemh("labels_10000.hex", all_labels);
        
        // �ʱ�ȭ
        rst_n = 0; valid_in = 0; data_in = 0;
        correct_cnt = 0;

        #100; rst_n = 1; #20;

        $display("\n========================================");
        $display(" Start Testing %0d Images...", NUM_TEST);
        $display("========================================\n");

        for (img_idx = 0; img_idx < NUM_TEST; img_idx = img_idx + 1) begin
            
            // �̹��� �ٲ� ������ ���� (�������� ���� ����)
            rst_n = 0; #20; rst_n = 1; #20;

            correct_label = all_labels[img_idx][3:0];
            base_addr = img_idx * 784;

            // �ȼ� ����
            for (px_idx = 0; px_idx < 784; px_idx = px_idx + 1) begin
                valid_in = 1;
                data_in = all_images[base_addr + px_idx];
                @(posedge clk); // ������ �������� ���� posedge ������ �ְ� ����ϰų�, ���⼭ ���
            end

            valid_in = 0;
            data_in = 0;

            // ��� ���
            wait(fc_done);
            @(posedge clk);

            // ä��
            if (final_digit == correct_label) begin
                correct_cnt = correct_cnt + 1;
            end else begin
                // Ʋ�� ��� �α� ��� (�ʹ� ���� ��µǸ� �ùķ��̼� �������Ƿ� �ʿ�� �ּ� ó��)
                // $display("Img %0d: FAIL (Pred: %d, True: %d)", img_idx, final_digit, correct_label);
            end
            
            // ���� ��Ȳ ��� (1000�� ������ ���� ��õ - 100���� �ʹ� ���� ����)
            if ((img_idx + 1) % 1000 == 0) begin
                $display("Process: %0d / %0d done... (Current Acc: %0.2f %%)", 
                         img_idx + 1, NUM_TEST, (correct_cnt * 100.0) / (img_idx + 1));
            end

            #200; // ���� �̹��� �� ������
        end

        $display("\n========================================");
        $display(" Test Finished!");
        $display(" Total Images: %0d", NUM_TEST);
        $display(" Correct     : %0d", correct_cnt);
        $display(" Accuracy    : %0.2f %%", (correct_cnt * 100.0) / NUM_TEST);
        $display("========================================");
        
        $finish;
    end

endmodule