module line_buffer_5x5 #(
    parameter DATA_BITS = 8,
    parameter WIDTH     = 28
)(
    input  wire                     clk,
    input  wire                     rst_n,
    input  wire [DATA_BITS-1:0]     data_in,
    input  wire                     data_valid,

    output reg  [DATA_BITS-1:0]     w00, w01, w02, w03, w04,
    output reg  [DATA_BITS-1:0]     w10, w11, w12, w13, w14,
    output reg  [DATA_BITS-1:0]     w20, w21, w22, w23, w24,
    output reg  [DATA_BITS-1:0]     w30, w31, w32, w33, w34,
    output reg  [DATA_BITS-1:0]     w40, w41, w42, w43, w44,

    output reg                      window_valid
);

    // ���� �޸�
    reg [DATA_BITS-1:0] line0 [0:WIDTH-1];
    reg [DATA_BITS-1:0] line1 [0:WIDTH-1];
    reg [DATA_BITS-1:0] line2 [0:WIDTH-1];
    reg [DATA_BITS-1:0] line3 [0:WIDTH-1];

    // ����Ʈ ��������
    reg [DATA_BITS-1:0] s0[0:4], s1[0:4], s2[0:4], s3[0:4], s4[0:4];

    integer i;
    reg [10:0] col_cnt; // �˳��ϰ� 11��Ʈ
    reg [10:0] row_cnt;

    always @(posedge clk or negedge rst_n) begin
      if (!rst_n) begin
        col_cnt <= 0;
        row_cnt <= 0;
        window_valid <= 0;
        // (�������� �ʱ�ȭ ���� ����, FPGA�� �ڵ� 0)
      end else if (data_valid) begin
        // 1. ������ �о�ֱ� (Shift)
        line3[col_cnt] <= line2[col_cnt];
        line2[col_cnt] <= line1[col_cnt];
        line1[col_cnt] <= line0[col_cnt];
        line0[col_cnt] <= data_in;

        for (i=4; i>0; i=i-1) begin
             s0[i] <= s0[i-1]; 
             s1[i] <= s1[i-1]; 
             s2[i] <= s2[i-1]; 
             s3[i] <= s3[i-1]; 
             s4[i] <= s4[i-1];
        end
        s0[0] <= data_in; 
        s1[0] <= line0[col_cnt]; 
        s2[0] <= line1[col_cnt]; 
        s3[0] <= line2[col_cnt]; 
        s4[0] <= line3[col_cnt];

        // 2. [����] �����ϰ� ���� ���� (������ ����)
        if (col_cnt == WIDTH-1) begin
            col_cnt <= 0;
            // �ٹٲ� �� ���� row ����
            if (row_cnt < 1000) row_cnt <= row_cnt + 1; 
        end else begin
            col_cnt <= col_cnt + 1;
        end

        // 3. ������ ��ȿ�� üũ (4�� �̻� �׿���, ���ε� 4ĭ �̻� ������ OK)
        // 3. �ڡڡ� [�ٽ� ����] ������ ��ȿ�� üũ (���� ����) �ڡڡ�
        // ����: 0~3��(4��)�� ä��� �� -> 4������ 27�������� ��ȿ
        // ����: 0~3��(4��)�� ä��� �� -> 4������ 27�������� ��ȿ
        if ((row_cnt >= 4 && row_cnt < WIDTH) && (col_cnt >= 4 && col_cnt < WIDTH))
            window_valid <= 1'b1;
        else
            window_valid <= 1'b0; // ���� ���̸� ��� ���� (Garbage Free)

      end else begin
        // �����Ͱ� �� ���� ���� valid�� ���ϴ� (���� ����)
        window_valid <= 1'b0; 
      end
    end

    // ��� ����
    always @(*) begin
        {w00,w01,w02,w03,w04} = {s4[4],s4[3],s4[2],s4[1],s4[0]};
        {w10,w11,w12,w13,w14} = {s3[4],s3[3],s3[2],s3[1],s3[0]};
        {w20,w21,w22,w23,w24} = {s2[4],s2[3],s2[2],s2[1],s2[0]};
        {w30,w31,w32,w33,w34} = {s1[4],s1[3],s1[2],s1[1],s1[0]};
        {w40,w41,w42,w43,w44} = {s0[4],s0[3],s0[2],s0[1],s0[0]};
    end

endmodule