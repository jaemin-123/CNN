`timescale 1ns / 1ps

module requantizer #(
    parameter IN_W = 32,
    parameter OUT_W = 8,
    parameter MULTIPLIER = 116,
    parameter SHIFT = 16
)(
    input wire clk,
    input wire rst_n,
    input wire valid_in,
    input wire signed [IN_W-1:0] data_in,
    output reg valid_out,
    output reg signed [OUT_W-1:0] data_out
);

    // ���� ����� ����Ʈ ����� ���� ����� ū �׸� (Overflow ����)
    reg signed [IN_W+15:0] scaled;  
    reg signed [IN_W+15:0] shifted; 

    // 8��Ʈ ���� (-128 ~ 127)
    localparam signed [IN_W+15:0] MAX_VAL = 127;
    localparam signed [IN_W+15:0] MIN_VAL = -128;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            valid_out <= 0;
            data_out <= 0;
            scaled <= 0;
            shifted <= 0;
        end else begin
            valid_out <= valid_in;
            
            if (valid_in) begin
                // 1. ���ϱ�
                scaled = data_in * $signed(MULTIPLIER);
                
                // 2. ������ (Arithmetic Shift: ��ȣ ����)
                shifted = scaled >>> SHIFT;
                
                // 3. �� �ٽ�: �ڸ��� ���� 32��Ʈ ���¿��� �˻� ��
                if (shifted > MAX_VAL) 
                    data_out <= 127;       // 127���� ũ�� 127�� ����
                else if (shifted < MIN_VAL) 
                    data_out <= -128;      // -128���� ������ -128�� ����
                else 
                    data_out <= shifted[OUT_W-1:0]; // ���� ���̸� ���� ��Ʈ�� ���
            end
        end
    end

endmodule