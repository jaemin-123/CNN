`timescale 1ns / 1ps

module parallel_to_serial #(
    parameter DATA_W = 8
)(
    input  wire clk,
    input  wire rst_n,
    
    // ���� �Է� (Layer 2�� ��� 3��)
    input  wire signed [DATA_W-1:0] din_0,
    input  wire signed [DATA_W-1:0] din_1,
    input  wire signed [DATA_W-1:0] din_2,
    input  wire vin_0, vin_1, vin_2, // �� ä���� Valid ��ȣ
    
    // ���� ��� (FC Layer�� ���� ��)
    output reg signed [DATA_W-1:0] dout,
    output reg vout
);

    reg signed [DATA_W-1:0] buf_1, buf_2; // ������ �ӽ� �����
    reg [1:0] state; // ���� ����� ���� ����

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= 0;
            vout  <= 0;
            dout  <= 0;
            buf_1 <= 0;
            buf_2 <= 0;
        end else begin
            vout <= 0; // �⺻������ 0 (Pulse)

            // 1. �� ���� ���ÿ� ������ ���� (Layer 2 �Ϸ� ����)
            if (vin_0 && vin_1 && vin_2) begin
                vout  <= 1;
                dout  <= din_0; // ù ��° ���� �ٷ� ������
                
                buf_1 <= din_1; // �� ��° �� ����
                buf_2 <= din_2; // �� ��° �� ����
                state <= 1;     // "������ �� ��° �� ���� ���ʾ�" ��� ���
            end 
            // 2. �����ص� �� ��° �� �߼�
            else if (state == 1) begin
                vout  <= 1;
                dout  <= buf_1;
                state <= 2;
            end
            // 3. �����ص� �� ��° �� �߼�
            else if (state == 2) begin
                vout  <= 1;
                dout  <= buf_2;
                state <= 0; // �ٽ� ��� ���·�
            end
        end
    end

endmodule