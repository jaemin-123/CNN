`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/12/22 11:50:09
// Design Name: 
// Module Name: fc
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fc_layer_digit_classifier (
    input clk,
    input valid_in,
    input signed [7:0] feature_in, // MaxPool���� ���� ������ �ϳ��� �Է�
    output reg [3:0] result_digit, // ���� �Ǻ��� ���� (0~9)
    output reg result_valid
);
    // 0~9�� Ŭ������ ���� ���� ������
    reg signed [31:0] scores [0:9];
    
    // ����ġ ROM (layer_3_weight)
    // �ּ�: {�Է� �ε���, Ŭ���� ��ȣ}
    wire signed [7:0] weight; 
    
    // ������ Ư¡ �����Ϳ� ���� ���� ��� (MAC ����)
    always @(posedge clk) begin
        if (valid_in) begin
            // ��� Ŭ����(0~9)�� ���� ���ÿ� ����ġ ���ؼ� ���ϱ�
            scores[0] <= scores[0] + feature_in * weight_0;
            scores[1] <= scores[1] + feature_in * weight_1;
            scores[2] <= scores[2] + feature_in * weight_2;
            scores[3] <= scores[3] + feature_in * weight_3;
            scores[4] <= scores[4] + feature_in * weight_4;
            scores[5] <= scores[5] + feature_in * weight_5;
            scores[6] <= scores[6] + feature_in * weight_6;
            scores[7] <= scores[7] + feature_in * weight_7;
            scores[8] <= scores[8] + feature_in * weight_8;
            scores[9] <= scores[9] + feature_in * weight_9;
        end
    end
    
    // ��� �Է��� ������ ���� ū ���� ã�� (ArgMax)
    always @(posedge clk) begin
        if (processing_done) begin
            // scores[0] ~ scores[9] �� �ִ밪�� �ε����� result_digit�� ����
        end
    end
endmodule
