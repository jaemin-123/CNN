`timescale 1ns / 1ps

module parallel_to_serial #(
    parameter DATA_W = 8
)(
    input  wire clk,
    input  wire rst_n,
    
    // ���� �Է�
    input  wire signed [DATA_W-1:0] din_0, din_1, din_2,
    input  wire vin_0, vin_1, vin_2, 
    
    // ���� ���
    output reg signed [DATA_W-1:0] dout, // reg ���� ���� (�����ϴ�!)
    output reg vout
);

    // 3���� ���� FIFO
    reg signed [DATA_W-1:0] q0 [0:63];
    reg signed [DATA_W-1:0] q1 [0:63];
    reg signed [DATA_W-1:0] q2 [0:63];

    reg [5:0] wp0, wp1, wp2; 
    reg [5:0] rp0, rp1, rp2; 
    
    // ������ ���� Ȯ�ο�
    wire [5:0] cnt0 = wp0 - rp0;
    wire [5:0] cnt1 = wp1 - rp1;
    wire [5:0] cnt2 = wp2 - rp2;

    reg [1:0] state; 

    // �ڡڡ� [����] Edge Detector ����! (�ܼ��ϰ� ���ϴ�) �ڡڡ�
    // reg vin_0_prev... ����
    // wire v0_pulse... ����

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            wp0 <= 0; wp1 <= 0; wp2 <= 0;
            rp0 <= 0; rp1 <= 0; rp2 <= 0;
            state <= 0;
            vout  <= 0;
            dout  <= 0;
            // vin_prev �ʱ�ȭ ����
        end else begin
            // 1. ���� (Pulse�� �ƴ϶� Valid�� ������ ����!)
            // �մ�(MaxPool)�� ��ȿ�� �����͸� �� �� �ϰ� �޽��ϴ�.
            if (vin_0) begin q0[wp0] <= din_0; wp0 <= wp0 + 1; end
            if (vin_1) begin q1[wp1] <= din_1; wp1 <= wp1 + 1; end
            if (vin_2) begin q2[wp2] <= din_2; wp2 <= wp2 + 1; end

            // 2. �б� (FSM - ������ ����)
            vout <= 0; 

            case (state)
                0: begin
                    // 3�� ä�� ��� �����Ͱ� 1�� �̻� ���� ���� ����
                    if (cnt0 > 0 && cnt1 > 0 && cnt2 > 0) begin
                        dout <= q0[rp0];     
                        vout <= 1;
                        rp0  <= rp0 + 1;     
                        state <= 1;          
                    end
                end
                
                1: begin
                    dout <= q1[rp1];        
                    vout <= 1;
                    rp1  <= rp1 + 1;        
                    state <= 2;             
                end

                2: begin
                    dout <= q2[rp2];        
                    vout <= 1;
                    rp2  <= rp2 + 1;        
                    state <= 0;             
                end
            endcase
        end
    end

endmodule