`timescale 1ns / 1ps

module preprocessing_unit (
    input  wire clk,
    input  wire rst_n,
    input  wire valid_in,
    input  wire [7:0] raw_data_in, // 0 ~ 255
    
    output reg  valid_out,
    output reg  signed [7:0] data_out // -19 ~ 127
);

    reg [15:0] mult_result;
    reg valid_stage1; // �� ���ڸ� ���߱� ���� �߰� Valid �������� �߰�

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            valid_stage1 <= 0;
            valid_out    <= 0;
            mult_result  <= 0;
            data_out     <= 0;
        end else begin
            // [Stage 1] ���� ����
            // valid_in ��ȣ�� ���� �� ���� ���� �� (valid_stage1�� ����)
            mult_result  <= raw_data_in * 147;
            valid_stage1 <= valid_in; 
            
            // [Stage 2] ���� ���� (���)
            // �����Ͱ� ���� �� valid_stage1�� valid_out���� ������ -> 2Ŭ�� �������� ��ũ ����
            data_out  <= mult_result[15:8] - 8'd19;
            valid_out <= valid_stage1; 
        end
    end

endmodule