`timescale 1ns / 1ps

module tb_latency_real();

    // 1. �Ķ���� �� ��ȣ ����
    reg clk;
    reg rst_n;
    reg valid_in;
    reg signed [7:0] data_in;
    
    wire fc_done;
    wire [3:0] final_digit;

    // 2. ������ ���� �� ���� ó�� ����
    real start_time;
    real end_time;
    real total_cycles;
    integer i;
    integer fd;         // ���� ��ũ����
    integer code;       // ���� �б� ����
    reg [7:0] pixel_temp; // ���Ͽ��� ���� �� �ӽ� ����

    // 3. DUT (Device Under Test) ����
    cnn_multichannel_top u_dut (
        .clk(clk),
        .rst_n(rst_n),
        .valid_in(valid_in),
        .data_in(data_in),
        .fc_done(fc_done),
        .final_digit(final_digit)
    );

    // 4. Ŭ�� ���� (125MHz = 8ns �ֱ�)
    always #4 clk = ~clk; 

    // 5. �׽�Ʈ �ó�����
    initial begin
        // �� [������ ����] ��� �Է� ��ȣ�� 0���� �ʱ�ȭ (���� �߿�)
        clk = 0;
        rst_n = 0;
        valid_in = 0;
        data_in = 0;
        pixel_temp = 0;

        // ���� ���� (Vivado ������Ʈ ���� -> simulation ���� �ȿ� ������ �־�� ��)
        fd = $fopen("raw_images_1000.hex", "r");
        if (fd == 0) begin
            $display("Error: 'raw_images_1000.hex' ������ ã�� �� �����ϴ�!");
            $stop;
        end

        // ���� ������ (����� �ð� ���� ���� ����)
        #100;
        rst_n = 1;
        #20;

        $display("========================================================");
        $display("[TB] Simulation Start: Measuring Inference Latency");
        $display("========================================================");

        // Ŭ�� ������ ���缭 ����
        @(posedge clk); 
        start_time = $time; // �� ���� �ð� ���

        // 6. ������ �Է� (���Ͽ��� ù ��° �̹��� 784 �ȼ��� ����)
        valid_in = 1;
        for (i = 0; i < 784; i = i + 1) begin
            // ��� ���Ͽ��� 1��(1�ȼ�) �б�
            code = $fscanf(fd, "%h", pixel_temp); 
            
            // ���� ������ �Է�
            data_in = pixel_temp;
            
            @(posedge clk);  // 1Ŭ�� ���
        end
        
        // �Է� ��
        valid_in = 0;
        data_in = 0;
        $fclose(fd); // ���� �ݱ�

        // 7. ��� ��� (fc_done�� 1�� �� ������)
        wait(fc_done == 1);
        
        // �� ���� �ð� ���
        end_time = $time; 

        // 8. ��� ��� �� ��� (���� ���� ����)
        // (����ð� - ���۽ð�) / Ŭ���ֱ�(8ns)
        total_cycles = (end_time - start_time) / 8.0;

        $display("========================================================");
        $display("[TB] Inference Completed!");
        $display("--------------------------------------------------------");
        $display("   - Start Time      : %0t ns", start_time);
        $display("   - End Time        : %0t ns", end_time);
        $display("   - Total Time      : %0t ns", (end_time - start_time));
        $display("--------------------------------------------------------");
        $display("�� Total Clock Cycles : %0d cycles", total_cycles);
        $display("========================================================");

        $stop; // �ùķ��̼� ����
    end

endmodule